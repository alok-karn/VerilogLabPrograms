module read_reg (
    clk, rst, ra, rb, busa, busb
);
    
endmodule